`ifndef F1_F2_PPREG
`define F1_F2_PPREG
    `include "f1_f2_ppreg.sv"
`endif