`ifndef FORWARDING_UNIT
`define FORWARDING_UNIT
    `include "internal_op.svh"
    `include "forwarding_unit.sv"
`endif