`ifndef SRAM_WRAPPER
`define SRAM_WRAPPER
    `include "SRAM_wrapper.sv"
    `include "SRAM_rtl.sv"
`endif