`ifndef D_E_PPREG
`define D_E_PPREG
    `include "d_e_ppreg.sv"
`endif