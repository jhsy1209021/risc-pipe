`ifndef MMU
`define MMU
    `include "mmu.sv"
    `include "internal_op.svh"
`endif