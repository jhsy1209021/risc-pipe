`ifndef BRANCH_COMPARATOR
`define BRANCH_COMPARATOR
    `include "branch_comparator.sv"
`endif