`ifndef F2_D_PPREG
`define F2_D_PPREG
    `include "f2_d_ppreg.sv"
`endif