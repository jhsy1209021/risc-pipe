`ifndef ALU
`define ALU
    `include "internal_op.svh"
`endif