`ifndef ALU
`define ALU
    `include "alu.sv"
    `include "internal_op.svh"
`endif