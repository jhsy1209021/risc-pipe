`ifndef CSR_ALU
`define CSR_ALU
    `include "internal_op.svh"
`endif
