`ifndef REGFILE
`define REGFILE
    `include "regfile.sv"
`endif