`ifndef ALU_OP
`define ALU_OP
    `define 
`endif