`ifndef FORWARDING_UNIT
`define FORWARDING_UNIT
    `include "forwarding_unit.sv"
    `include "internal_op.svh"
`endif