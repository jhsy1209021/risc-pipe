`ifndef E_M1_PPREG
`define E_M1_PPREG
    `include "e_m1_ppreg.sv"
`endif