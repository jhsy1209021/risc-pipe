`ifndef READ_ALIGNER
`define READ_ALIGNER
    `include "internal_op.svh"
    `include "read_aligner.sv"
`endif