`ifndef HAZARD_ELIMINATOR
`define HAZARD_ELIMINATOR
    `include "internal_op.svh"
    `include "hazard_eliminator.sv"
`endif