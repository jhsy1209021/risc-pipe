`ifndef SRAM_WRAPPER
`define SRAM_WRAPPER
    `include "SRAM_rtl.sv"
    `include "SRAM_wrapper.sv"
`endif