`ifndef HAZARD_ELEMINATOR
`define HAZARD_ELEMINATOR
    `include "hazard_eleiminator.sv"
    `include "internal_op.svh"
`endif