`ifndef ALU
`define ALU
    `include "internal_op.svh"
    `include "alu.sv"
`endif