`ifndef WB_UNIT
`define WB_UNIT
    `include "wb_unit.sv"
    `include "internal_op.svh"
`endif