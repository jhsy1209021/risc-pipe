`ifndef SRAM_WRAPPER
`define SRAM_WRAPPER
    `include "SRAM_wrapper.sv"
`endif