`ifndef ADDR_GEN
`define ADDR_GEN
    `include "addr_gen.sv"
`endif