`ifndef MMU
`define MMU
    `include "internal_op.svh"
`endif