`ifndef M2_WB_PPREG
`define M2_WB_PPREG
    `include "m2_wb_ppreg.sv"
`endif