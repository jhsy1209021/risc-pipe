`ifndef CSR_REG_BANK
`define CSR_REG_BANK
    `include "csr_reg_bank.sv"
`endif