`ifndef PC
`define PC
    `include "pc.sv"
`endif