`ifndef READ_ALIGNER
`define READ_ALIGNER
    `include "read_aligner.sv"
    `include "internal_op.svh"
`endif