`ifndef HAZARD_ELIMINATOR
`define HAZARD_ELIMINATOR
    `include "hazard_eliminator.sv"
    `include "internal_op.svh"
`endif