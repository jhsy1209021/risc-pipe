`ifndef WB_UNIT
`define WB_UNIT
    `include "internal_op.svh"
    `include "wb_unit.sv"
`endif