`ifndef CSR_ALU
`define CSR_ALU
    `include "csr_alu.sv"
    `include "internal_op.svh"
`endif
