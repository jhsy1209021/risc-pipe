`ifndef MMU
`define MMU
    `include "internal_op.svh"
    `include "mmu.sv"
`endif