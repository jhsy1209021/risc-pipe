`ifndef M1_M2_PPREG
`define M1_M2_PPREG
    `include "m1_m2_ppreg.sv"
`endif